
* Project HARLEMSHAKEDETECTOR
* Mentor Graphics Netlist Created with Version 5.8
* File created Mon Mar 11 14:59:28 2013
* Inifile   : 
*
* Config file: C:\MentorGraphics\SystemVision5.9\standard\svspice.cfg
*
* Options   : -_ -h -kC:\MentorGraphics\SystemVision5.9\standard\svspice.cfg -gharlemshakedetector.tempfile 
* 
* Levels    : 
* 
.option noinclib
* Models for Eldo<->VHDL-AMS data conversion
.model a2d_eldo a2d mode=std_logic VTH=1.65
.model d2a_eldo d2a mode=std_logic VHI=3.3 VLO=0.0
.defhook a2d_eldo
.defhook d2a_eldo
.param process_corner=0
YV3 V_CONSTANT(IDEAL) GENERIC: LEVEL="1.65" PORT: AVDD VCM
YAL1 VIA_DL_DFFR(LEVEL_2) GENERIC: DELAY="0.1800E-9" SIGNALTYPE="ANALOG" PORT: 
+ AVDD DEEP_VOICE_DETECTED AVDD DO_THE_HARLEM_SHAKE
YN1I43 V_VS_TIME_FROM_FILE(IDEAL) PORT: MUSIC VCM
YV1 V_CONSTANT(IDEAL) GENERIC: LEVEL="0.0" PORT: AVSS 0
YFLTR2 VIA_FILTER_CONTINUOUS(LEVEL_0) GENERIC: 
+ A="(8.76995679608E+59,7.62397855445E+56,1.18475482273E+55,9.10242494647E+51,6.82744365675E+49,4.56165284385E+46,2.1957548253E+44,1.25002687542E+41,4.33682265797E+38,2.04996861625E+35,5.46958267798E+32,2.07705246628E+29,4.45217444485E+26,1.3002297964E+23,2.31411461013E+20,4.87106028026E+16,7.3868563328E+13,9978353579.54,13159231.3467,857.993420542,1.0)" 
+ AREA="3070200" 
+ B="(8.76688554048E+56,0.0,2.49811726295E+52,0.0,2.40350009005E+47,0.0,1.11661512337E+42,0.0,2.79493536401E+36,0.0,3.84917080404E+30,0.0,2.869275685E+24,0.0,1.17680505179E+18,0.0,260043301032.0,0.0,27746.9248182,0.0,0.000999649798092)" 
+ BW="150.0" FC="158.1" FILTERTYPE="BANDPASS" FSTOP="250" ISUPNOM="9500" 
+ ORDER="10" SETTLETIME="(5.6E-06,1E-06,1E-05)" STOPATTEN="60" STYLE="ELLIP" 
+ PORT: AVDD MUSIC DEEP_VOICE_FILTERED AVDD AVSS VCM
YCMP1 VIA_CMP_OA(LEVEL_0) GENERIC: GM="(12.7E-3,10.8E-3,14.86E-3)" VHYST="50" 
+ PORT: AVDD AVSS DEEP_VOICE_DETECTED AVDD SLICE_LEVEL DEEP_VOICE_FILTERED
YV4 V_CONSTANT(IDEAL) GENERIC: LEVEL="1.7" PORT: SLICE_LEVEL 0
YV2 V_CONSTANT(IDEAL) GENERIC: LEVEL="1.65" PORT: VCM AVSS
* DICTIONARY 1
* GND = 0
*Note: Floating node DO_THE_HARLEM_SHAKE.
.GLOBAL ELECTRICAL_REF
.model V_VS_TIME_FROM_FILE(IDEAL) macro lang=vhdlams LIB=EDULIB
.model V_CONSTANT(IDEAL) macro lang=vhdlams LIB=EDULIB
.model VIA_FILTER_CONTINUOUS(LEVEL_0) macro lang=vhdlams LIB=WORK
.model VIA_CMP_OA(LEVEL_0) macro lang=vhdlams LIB=WORK
.model VIA_DL_DFFR(LEVEL_2) macro lang=vhdlams LIB=WORK
.END
